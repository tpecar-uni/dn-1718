`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:52:23 02/06/2017 
// Design Name: 
// Module Name:    dataSyncModule 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module dataSyncModule(
    input clk_i,
    input reset_i,
    input clksync_i,
    output pulse_o
    );


endmodule
